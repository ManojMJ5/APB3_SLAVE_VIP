package apb_pkg;
`include "uvm_macros.svh"
 import uvm_pkg::*;

`include "apb_seqitems.sv"
`include "apb_sequence.sv"
`include "apb_sequencer.sv"
`include "apb_driver.sv"
`include "apb_imonitor.sv"
`include "apb_iagent.sv"
`include "apb_sb_predictor.sv"
`include "apb_sb_comparator.sv"
`include "apb_scoreboard.sv"
`include "apb_coverage.sv"
`include "apb_env.sv"
`include "base_test.sv"
endpackage
