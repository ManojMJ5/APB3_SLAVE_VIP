`define CYCLE 10
`define TDRIVE #(0.8 * `CYCLE)
`timescale 1ns/1ns